module rx_fifo(

);




endmodule