module rxfifo_tb();





endmodule